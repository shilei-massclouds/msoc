`timescale 1ns / 1ps

`include "isa.vh"

module regfile (
    input  wire         clk,
    input  wire         rst_n,

    input  wire [4:0]   rs1,
    output wire [63:0]  data1,
    input  wire [4:0]   rs2,
    output wire [63:0]  data2,
    input  wire [4:0]   wb_rd,
    input  wire [63:0]  wb_data
);

    reg [63:0] data[32];

    assign data1 = (rs1 == 5'b0) ? 64'b0 :
                   (rs1 == wb_rd) ? wb_data : data[rs1];

    assign data2 = (rs2 == 5'b0) ? 64'b0 :
                   (rs2 == wb_rd) ? wb_data : data[rs2];

    always @(posedge clk, negedge rst_n) begin
        if (~rst_n) begin
            for (integer i = 0; i < 32; i++)
                data[i] <= 64'b0;
        end else begin
            if (wb_rd) data[wb_rd] <= wb_data;
        end
    end

endmodule
